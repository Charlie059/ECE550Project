/* This module is a NOT GATE
Xuhui Gong	21-09-11
*/
module NOT_1(out, in);
	
	input in;
	output out;
	
	not not_gate(out, in);

endmodule